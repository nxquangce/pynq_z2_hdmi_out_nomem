`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Computer Engineering Lab - CSE - HCMUT
// Engineer: Nguyen Xuan Quang
// 
// Create Date: 11/24/2020 11:15:15 AM
// Design Name: pynq-z2-hdmi-out-nomem
// Module Name: top
// Project Name: pynq-z2-hdmi-out-nomem
// Target Devices: pynq-x2
// Tool Versions: 2018.2
// Description: pynq-z2-hdmi-out-nomem top module
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(
    DDR_addr,
    DDR_ba,
    DDR_cas_n,
    DDR_ck_n,
    DDR_ck_p,
    DDR_cke,
    DDR_cs_n,
    DDR_dm,
    DDR_dq,
    DDR_dqs_n,
    DDR_dqs_p,
    DDR_odt,
    DDR_ras_n,
    DDR_reset_n,
    DDR_we_n,
    FIXED_IO_ddr_vrn,
    FIXED_IO_ddr_vrp,
    FIXED_IO_mio,
    FIXED_IO_ps_clk,
    FIXED_IO_ps_porb,
    FIXED_IO_ps_srstb,
    TMDS_Clk_n_0,
    TMDS_Clk_p_0,
    TMDS_Data_n_0,
    TMDS_Data_p_0,
    led
);

    parameter DATA_WIDTH     = 24;
    parameter ROW_ADDR_WIDTH = 10;
    parameter COL_ADDR_WIDTH = 11;
    parameter PATTERN_MODE   = 1;
    parameter MAX_COL        = 1280;   // 800, 1280
    parameter MAX_ROW        = 1024;   // 600, 1024

    inout [14:0]    DDR_addr;
    inout [2:0]     DDR_ba;
    inout           DDR_cas_n;
    inout           DDR_ck_n;
    inout           DDR_ck_p;
    inout           DDR_cke;
    inout           DDR_cs_n;
    inout [3:0]     DDR_dm;
    inout [31:0]    DDR_dq;
    inout [3:0]     DDR_dqs_n;
    inout [3:0]     DDR_dqs_p;
    inout           DDR_odt;
    inout           DDR_ras_n;
    inout           DDR_reset_n;
    inout           DDR_we_n;
    inout           FIXED_IO_ddr_vrn;
    inout           FIXED_IO_ddr_vrp;
    inout [53:0]    FIXED_IO_mio;
    inout           FIXED_IO_ps_clk;
    inout           FIXED_IO_ps_porb;
    inout           FIXED_IO_ps_srstb;
    output          TMDS_Clk_n_0;
    output          TMDS_Clk_p_0;
    output [2:0]    TMDS_Data_n_0;
    output [2:0]    TMDS_Data_p_0;
    output [3:0]    led;

    wire [14:0]     DDR_addr;
    wire [2:0]      DDR_ba;
    wire            DDR_cas_n;
    wire            DDR_ck_n;
    wire            DDR_ck_p;
    wire            DDR_cke;
    wire            DDR_cs_n;
    wire [3:0]      DDR_dm;
    wire [31:0]     DDR_dq;
    wire [3:0]      DDR_dqs_n;
    wire [3:0]      DDR_dqs_p;
    wire            DDR_odt;
    wire            DDR_ras_n;
    wire            DDR_reset_n;
    wire            DDR_we_n;
    wire            FIXED_IO_ddr_vrn;
    wire            FIXED_IO_ddr_vrp;
    wire [53:0]     FIXED_IO_mio;
    wire            FIXED_IO_ps_clk;
    wire            FIXED_IO_ps_porb;
    wire            FIXED_IO_ps_srstb;
    wire            TMDS_Clk_n_0;
    wire            TMDS_Clk_p_0;
    wire [2:0]      TMDS_Data_n_0;
    wire [2:0]      TMDS_Data_p_0;
    wire [3:0]      led;
  
    wire                      clk_100M;
    wire [ROW_ADDR_WIDTH-1:0] row_address;
    wire [COL_ADDR_WIDTH-1:0] col_address;
    wire [DATA_WIDTH-1:0]     video_data;
    wire                      next_pixel;

    video_out_pynq_z2_wrapper video_out_pynq_z2_wrapper_i (
        .DDR_addr           (DDR_addr),
        .DDR_ba             (DDR_ba),
        .DDR_cas_n          (DDR_cas_n),
        .DDR_ck_n           (DDR_ck_n),
        .DDR_ck_p           (DDR_ck_p),
        .DDR_cke            (DDR_cke),
        .DDR_cs_n           (DDR_cs_n),
        .DDR_dm             (DDR_dm),
        .DDR_dq             (DDR_dq),
        .DDR_dqs_n          (DDR_dqs_n),
        .DDR_dqs_p          (DDR_dqs_p),
        .DDR_odt            (DDR_odt),
        .DDR_ras_n          (DDR_ras_n),
        .DDR_reset_n        (DDR_reset_n),
        .DDR_we_n           (DDR_we_n),
        .FIXED_IO_ddr_vrn   (FIXED_IO_ddr_vrn),
        .FIXED_IO_ddr_vrp   (FIXED_IO_ddr_vrp),
        .FIXED_IO_mio       (FIXED_IO_mio),
        .FIXED_IO_ps_clk    (FIXED_IO_ps_clk),
        .FIXED_IO_ps_porb   (FIXED_IO_ps_porb),
        .FIXED_IO_ps_srstb  (FIXED_IO_ps_srstb),
        .TMDS_Clk_n_0       (TMDS_Clk_n_0),
        .TMDS_Clk_p_0       (TMDS_Clk_p_0),
        .TMDS_Data_n_0      (TMDS_Data_n_0),
        .TMDS_Data_p_0      (TMDS_Data_p_0),

        // User port
        .clk_100M           (clk_100M),
        .col_address        (col_address),
        .data_in            (video_data),
        .next_pixel         (next_pixel),
        .row_address        (row_address)
    );

    video_pattern_generator
    #(
        .DATA_WIDTH     (DATA_WIDTH),
        .ROW_ADDR_WIDTH (ROW_ADDR_WIDTH),
        .COL_ADDR_WIDTH (COL_ADDR_WIDTH),
        .PATTERN_MODE   (PATTERN_MODE),
        .MAX_ROW        (MAX_ROW),
        .MAX_COL        (MAX_COL)
    )
    video_pattern_generator_i
    (
        .clk            (clk_100M),
        .next_pixel     (next_pixel),
        .row_address    (row_address),
        .col_address    (col_address),
        .data_out       (video_data)
    );
endmodule
